module dut2 (
    input a,
    output b
);

assign b = ~a;

endmodule
